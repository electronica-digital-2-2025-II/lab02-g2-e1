`include "four_adder.v"
`include "adder.v"
`include "mult.v"
`include "shift.v"

module alu(
    input clk,
    input [3:0] a,
    input [3:0] b,
    input [2:0] op,
    input init,
    input cin,
    
    output reg [6:0] result,
    output reg carry,
    output reg done,
    output reg overflow,
    output reg zero
);

    wire done_;
    wire carry_;
    wire [3:0] sum_;
    wire [6:0] sum_result = {carry_, sum_};
    wire [7:0] mul_result;
    wire [6:0] shift_w;
    wire [6:0] rest_result = {2'b00, sum_};
    reg [6:0] temp_result;

    // Instancias
    four_adder sum(
        .a(a),
        .b(b),
        .cin(cin),
        .sum(sum_),
        .carry(carry_)
    );

    shift sh(
        .a(a),
        .shift_(b),
        .shift_number(shift_w),
        .done(done_)
    );

    mult mul(
        .a(a),
        .b(b),
        .clk(clk),
        .init(init),
        .result(mul_result),
        .done(done_)
    );

    always @(posedge clk) begin
        
        if (init) begin
            result <= 7'b0000000;
            overflow <= 1'b0;
            done <= 1'b0;
            carry <= 1'b0;
            zero <= 1'b0;

        end else begin
            temp_result = 7'b0000000;
            overflow = 1'b0;
            carry = 1'b0;
            done = 1'b0;

            case (op)
                3'b001: begin // Suma
                    if (cin) begin
                        temp_result = rest_result;
                        carry = carry_;

                    end else begin
                        temp_result = sum_result;
                        carry = carry_;
                    end
                end

                3'b010: begin // Multiplicación
                    temp_result = mul_result[6:0];
                    overflow = mul_result[7];
                    done = done_;
                end

                3'b011: begin // Desplazamiento
                    temp_result = shift_w;
                    done = done_;
                end

                3'b111: begin // Operación lógica: AND
                    temp_result = a & b;
                    done = done_;
                end

                default: begin
                    temp_result = 7'b0000000;
                    overflow = 1'b0;
                end
            endcase

            // Salidas 
            result <= temp_result;
            zero <= (temp_result == 0);
            carry <= carry;
            overflow <= overflow;
            done <= done;
        end
    end

endmodule